enum bit [6:0] {
  AND  = 0, 
  ANDN = 1, 
  OR   = 2, 
  ORN  = 3, 
  XOR  = 4, 
  XORN = 5, 
  NOT  = 6, 
  ADD  = 7, 
  SUB  = 8, 
  MUL  = 9, 
  DIV  = 10, 
  MOD  = 11, 
  GT   = 12, 
  GE   = 13, 
  EQ   = 14, 
  NE   = 15, 
  LE   = 16, 
  LT   = 17, 
  JMP  = 18, 
  IF0JUMP = 19,     
  IF1JUMP = 20,     
  CALL  = 21,      
  CAL0 = 22, 
  CAL1 = 23, 
  RET  = 24,       
  RET0 = 25,
  RET1 = 26,
  SET = 27,
  RST = 28,      
  ST = 29,
  STN = 30,
  LD = 31,
  LDN = 32
}opCodes;
