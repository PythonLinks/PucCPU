   initial
     $monitor ("%f", position,  " ",
	        velocity , " ",
           scaledPosition, " ",
	       positionOutInt, " ",
               positionOut);
