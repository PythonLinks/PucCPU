`ifndef GLOBAL
//`define DEMO1 1
//`define DEMO2 1
`define PBL 1
`define GLOBAL 1
`endif  
